LIBRARY ieee;
USE work.twoD_array.ALL;

ENTITY filter_tb IS
END filter_tb;

ARCHITECTURE test OF filter_tb IS
	COMPONENT sharp_filter IS
		GENERIC(n : INTEGER := 32;
				m : INTEGER := 64);
		PORT(
			input    : IN  array_2d(0 TO n-1,0 TO m-1);
			output_1 : OUT array_2d(0 TO n-1,0 TO m-1);
		    output_2 : OUT array_2d(0 TO n-1,0 TO m-1)		
		);	
	END COMPONENT;
	
SIGNAL input_t : array_2d(0 TO 31,0 TO 63) := ((130,130,130,131,131,130,132,132,131,122,89,54,16,3,2,1,2,2,7,36,69,96,104,105,106,106,107,108,109,109,110,109,110,112,103,35,10,11,11,13,37,64,66,66,66,67,68,67,67,68,66,68,68,68,69,40,14,12,10,10,10,10,9,11),
(130,130,131,132,131,132,132,132,133,133,132,131,58,2,1,2,3,3,44,100,104,104,104,104,106,107,107,107,110,108,111,110,110,99,32,11,11,10,12,25,63,66,65,66,66,65,66,67,67,68,68,67,67,68,69,65,21,12,11,10,11,10,10,11),
(129,131,131,132,130,132,132,133,133,133,132,97,8,3,3,4,3,18,92,103,103,104,105,105,105,106,107,107,109,108,109,110,86,24,9,10,10,11,19,56,64,65,66,65,67,66,65,65,66,66,67,68,67,68,68,69,50,12,11,11,11,9,10,10),
(129,130,129,130,131,131,133,133,132,133,123,29,4,4,3,2,8,66,103,104,104,105,104,105,106,107,107,107,108,108,102,58,14,9,9,10,11,16,54,65,65,66,66,65,68,66,66,67,66,67,68,68,67,68,69,70,67,27,11,10,10,10,11,10),
(128,129,130,130,130,131,130,132,133,130,60,6,4,4,4,4,37,100,102,105,104,104,104,106,106,105,106,108,105,75,25,10,10,10,9,11,18,52,65,66,65,65,67,65,66,66,67,65,66,67,66,67,67,69,70,69,69,57,14,11,10,10,9,11),
(129,128,129,130,130,131,131,132,132,94,10,5,4,3,4,16,89,103,102,103,104,104,103,105,104,104,102,71,30,10,9,8,10,10,11,23,56,65,64,65,66,65,65,66,66,66,67,67,66,67,66,67,67,68,67,68,68,67,31,12,9,11,10,10),
(104,123,129,129,131,131,131,131,115,23,6,5,4,4,6,66,102,102,102,104,104,105,104,101,81,51,17,10,8,8,9,8,10,13,34,60,63,65,65,65,65,65,66,65,65,67,67,66,67,66,68,68,68,67,68,68,68,69,56,14,12,11,10,9),
(8,13,33,57,78,97,113,121,43,6,5,5,4,4,39,100,102,103,101,99,87,67,43,18,8,8,8,7,9,9,9,10,19,48,62,61,62,64,65,65,66,65,65,65,66,66,65,66,66,67,67,66,67,68,67,68,68,68,68,27,11,11,12,11),
(6,6,4,6,7,7,9,10,6,5,3,4,5,10,67,70,60,45,30,14,8,7,7,8,8,9,8,10,9,10,17,40,59,63,60,62,63,64,63,65,66,66,66,65,65,66,67,66,67,66,65,66,68,68,68,68,68,68,68,46,11,11,11,10),
(4,5,6,6,5,5,5,5,5,6,4,5,4,6,7,6,6,6,8,6,7,6,7,7,8,8,9,11,21,41,59,61,63,62,65,64,63,62,64,64,64,64,65,66,65,65,66,65,66,66,65,67,65,67,68,67,67,69,68,60,14,12,11,12),
(6,5,6,5,4,5,6,5,4,5,5,5,5,5,5,6,7,5,7,8,8,7,7,8,9,16,32,51,63,78,96,108,116,119,118,113,103,85,71,68,65,65,66,66,66,66,64,64,66,66,67,65,68,66,68,68,67,68,68,68,19,11,11,11),
(8,7,6,5,7,5,5,5,4,5,7,6,5,5,6,6,6,8,7,8,9,13,21,34,48,63,89,121,147,156,159,158,158,159,159,160,160,159,157,137,108,77,66,65,65,65,66,64,66,65,65,66,66,67,66,68,67,67,69,70,25,13,12,12),
(110,83,59,35,15,6,5,6,5,6,6,8,6,8,10,12,17,23,30,38,47,56,59,65,96,140,156,157,157,157,156,150,140,136,137,144,153,159,161,160,161,159,127,83,67,67,66,65,64,66,65,65,65,66,66,65,66,67,67,67,25,13,12,12),
(137,137,137,135,91,11,5,7,6,21,44,45,47,50,53,54,56,56,56,58,57,59,83,136,155,155,156,151,124,98,75,63,63,63,64,65,67,80,104,136,159,161,161,159,121,72,66,65,65,65,65,67,65,66,67,67,66,66,65,65,20,12,12,12),
(137,137,122,60,11,7,7,7,18,50,53,55,56,54,54,55,55,57,56,59,63,109,151,154,155,145,105,71,63,63,61,61,63,63,61,62,63,63,63,65,79,122,157,162,163,149,90,66,66,65,65,66,65,63,64,65,65,68,67,60,14,11,12,12),
(102,63,19,8,8,7,7,21,48,53,55,55,53,56,56,56,56,57,58,67,124,152,154,150,112,68,62,62,60,60,61,62,63,62,63,62,63,63,64,64,63,65,81,135,162,162,159,105,67,65,65,65,66,64,66,67,65,67,66,44,13,12,12,14),
(9,8,9,8,9,8,27,50,53,54,55,56,52,55,55,55,58,58,64,126,152,153,137,81,60,61,61,61,60,61,61,66,65,66,65,66,65,64,63,64,63,66,65,66,109,158,161,160,112,68,66,65,67,64,65,66,67,67,52,17,12,12,13,13),
(9,8,8,9,14,37,51,52,52,54,55,54,53,55,54,56,56,62,121,152,152,124,69,60,60,58,60,59,62,61,64,144,153,152,152,150,149,122,64,63,62,65,64,64,66,92,153,161,160,110,65,64,63,65,66,65,67,54,17,14,13,13,14,15),
(9,9,14,32,48,53,52,52,52,53,54,55,54,55,56,56,59,105,149,150,117,64,59,60,59,59,60,60,60,61,66,146,156,156,156,157,158,133,65,62,64,63,64,64,63,66,88,153,161,157,98,66,64,63,65,66,65,30,13,13,12,13,15,35),
(12,9,30,54,52,51,53,53,54,55,54,55,55,55,56,58,81,145,150,117,63,59,60,60,59,59,58,61,61,61,64,146,155,155,156,157,157,136,65,62,64,63,63,63,65,65,64,90,157,160,153,80,64,64,66,65,65,27,13,13,14,14,45,156),
(14,11,40,53,52,52,53,54,53,53,54,53,55,54,56,62,129,148,147,121,116,109,108,104,100,98,95,91,86,84,83,147,155,156,156,156,157,139,71,67,67,67,67,66,67,65,66,66,105,159,159,134,67,65,65,64,64,26,12,14,15,15,124,119),
(12,12,47,52,52,54,52,53,52,54,54,53,54,54,55,91,145,146,147,147,149,149,149,149,150,151,150,151,152,153,153,153,155,154,155,156,156,156,153,153,153,152,149,149,147,145,143,140,139,157,160,158,101,64,63,64,66,26,14,14,12,16,43,19),
(12,17,50,51,50,50,52,51,51,52,52,54,53,55,60,128,145,129,113,117,121,122,127,128,133,135,138,141,143,146,148,150,150,152,154,154,156,155,156,156,157,157,157,158,157,158,158,159,159,158,159,159,145,68,65,65,64,25,13,14,13,16,116,89),
(11,21,50,49,51,51,51,52,52,52,53,54,54,55,81,143,142,74,58,57,58,57,59,57,57,59,59,61,61,61,63,65,66,67,71,73,75,79,81,85,89,92,94,97,99,102,105,108,110,114,135,158,159,99,65,64,64,25,14,14,14,18,149,174),
(12,27,50,52,50,51,52,53,52,51,52,54,55,55,110,143,121,58,56,55,55,57,58,58,58,59,58,58,59,59,59,60,58,61,62,62,61,62,63,63,62,63,62,64,62,64,63,63,64,64,76,152,158,137,66,64,63,25,14,14,15,18,150,174),
(11,31,51,51,50,50,51,52,52,53,53,54,55,60,133,144,97,58,56,56,55,56,57,56,58,58,57,58,57,59,59,59,60,60,60,61,62,61,62,61,61,62,61,61,62,62,62,63,64,63,63,116,158,156,79,63,62,25,15,15,14,17,124,109),
(12,36,50,50,50,50,51,52,52,52,52,53,55,74,142,141,76,56,57,56,56,55,56,56,57,58,58,58,58,59,58,58,60,60,61,60,58,61,61,60,61,62,61,61,62,62,63,61,64,61,62,81,155,157,105,63,63,24,16,13,14,18,40,22),
(12,39,49,50,51,49,51,52,51,52,53,54,54,90,142,137,64,57,57,57,57,56,56,56,57,58,57,58,58,58,58,59,59,59,60,59,60,60,60,62,61,62,62,62,63,63,63,61,61,62,64,65,140,156,128,63,62,25,15,14,14,18,122,101),
(12,40,50,50,50,50,50,51,51,52,54,54,55,101,141,134,85,80,77,74,71,69,64,64,62,61,61,59,60,60,60,60,59,60,58,59,59,61,61,62,62,63,62,63,62,62,62,63,61,62,62,63,118,157,145,66,63,25,14,13,14,18,151,171),
(14,42,49,49,48,50,50,52,51,51,52,54,56,108,141,142,142,142,143,143,144,144,144,143,143,140,139,135,132,129,125,69,58,59,58,59,59,62,109,121,118,116,115,112,111,108,105,103,100,99,96,94,121,156,152,72,63,23,14,14,15,18,152,170),
(15,42,51,50,51,51,50,51,51,52,53,52,55,113,140,142,142,142,142,143,144,144,144,145,146,146,146,147,148,148,147,77,58,58,59,60,59,62,130,151,152,153,153,154,153,154,154,154,154,154,153,154,155,156,155,80,62,22,14,13,15,18,114,94),
(206,0,0,206,51,50,51,51,52,51,50,53,54,115,139,141,141,142,141,143,143,144,144,146,145,146,146,146,148,147,147,79,58,58,59,58,59,62,130,151,152,152,151,153,153,152,153,154,153,153,153,153,154,155,154,86,61,23,14,14,14,18,37,19));
SIGNAL output_1_t : array_2d(0 TO 31,0 TO 63);
SIGNAL output_2_t : array_2d(0 TO 31,0 TO 63);
	
BEGIN
lab: sharp_filter GENERIC MAP(32,64) PORT MAP (input_t,output_1_t,output_2_t);	
	
END test;
